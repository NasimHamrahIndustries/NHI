`timescale 1 ns/100 ps
// Version: v11.8 SP3 11.8.3.6


module FIFOCore_2Bto1B_2048(
       DATA,
       Q,
       WE,
       RE,
       CLK,
       FULL,
       EMPTY,
       RESET
    );
input  [15:0] DATA;
output [7:0] Q;
input  WE;
input  RE;
input  CLK;
output FULL;
output EMPTY;
input  RESET;

    wire READ_RESET_P, \MEM_RADDR[0] , \MEM_RADDR[1] , \MEM_RADDR[2] , 
        \MEM_RADDR[3] , \MEM_RADDR[4] , \MEM_RADDR[5] , \MEM_RADDR[6] , 
        \MEM_RADDR[7] , \MEM_RADDR[8] , \MEM_RADDR[9] , 
        \MEM_RADDR[10] , \MEM_RADDR[11] , \MEM_RADDR[12] , 
        \RBINNXTSHIFT[0] , \RBINNXTSHIFT[1] , \RBINNXTSHIFT[2] , 
        \RBINNXTSHIFT[3] , \RBINNXTSHIFT[4] , \RBINNXTSHIFT[5] , 
        \RBINNXTSHIFT[6] , \RBINNXTSHIFT[7] , \RBINNXTSHIFT[8] , 
        \RBINNXTSHIFT[9] , \RBINNXTSHIFT[10] , \RBINNXTSHIFT[11] , 
        \RBINNXTSHIFT[12] , \WBINSYNCSHIFT[1] , \WBINSYNCSHIFT[2] , 
        \WBINSYNCSHIFT[3] , \WBINSYNCSHIFT[4] , \WBINSYNCSHIFT[5] , 
        \WBINSYNCSHIFT[6] , \WBINSYNCSHIFT[7] , \WBINSYNCSHIFT[8] , 
        \WBINSYNCSHIFT[9] , \WBINSYNCSHIFT[10] , \WBINSYNCSHIFT[11] , 
        \WBINSYNCSHIFT[12] , \WBINNXTSHIFT[0] , \WBINNXTSHIFT[1] , 
        \WBINNXTSHIFT[2] , \WBINNXTSHIFT[3] , \WBINNXTSHIFT[4] , 
        \WBINNXTSHIFT[5] , \WBINNXTSHIFT[6] , \WBINNXTSHIFT[7] , 
        \WBINNXTSHIFT[8] , \WBINNXTSHIFT[9] , \WBINNXTSHIFT[10] , 
        \WBINNXTSHIFT[11] , FULLINT, MEMORYWE, MEMWENEG, \WGRY[0] , 
        \WGRY[1] , \WGRY[2] , \WGRY[3] , \WGRY[4] , \WGRY[5] , 
        \WGRY[6] , \WGRY[7] , \WGRY[8] , \WGRY[9] , \WGRY[10] , 
        \WGRY[11] , EMPTYINT, MEMORYRE, MEMRENEG, DVLDI, DVLDX, 
        \RGRY[0] , \RGRY[1] , \RGRY[2] , \RGRY[3] , \RGRY[4] , 
        \RGRY[5] , \RGRY[6] , \RGRY[7] , \RGRY[8] , \RGRY[9] , 
        \RGRY[10] , \RGRY[11] , \RGRY[12] , \QXI[0] , \QXI[1] , 
        \QXI[2] , \QXI[3] , \QXI[4] , \QXI[5] , \QXI[6] , \QXI[7] , 
        XOR2_11_Y, XOR2_20_Y, XOR2_40_Y, XOR2_41_Y, XOR2_59_Y, 
        XOR2_67_Y, XOR2_51_Y, XOR2_16_Y, XOR2_50_Y, XOR2_29_Y, 
        XOR2_62_Y, XOR2_4_Y, XOR2_30_Y, AND2_33_Y, AND2_16_Y, 
        AND2_43_Y, AND2_4_Y, AND2_15_Y, AND2_1_Y, AND2_28_Y, AND2_22_Y, 
        AND2_31_Y, AND2_24_Y, AND2_30_Y, AND2_54_Y, XOR2_53_Y, 
        XOR2_5_Y, XOR2_9_Y, XOR2_2_Y, XOR2_10_Y, XOR2_23_Y, XOR2_48_Y, 
        XOR2_3_Y, XOR2_12_Y, XOR2_60_Y, XOR2_46_Y, XOR2_6_Y, XOR2_68_Y, 
        AND2_17_Y, AO1_29_Y, AND2_50_Y, AO1_8_Y, AND2_18_Y, AO1_36_Y, 
        AND2_29_Y, AO1_31_Y, AND2_45_Y, AO1_15_Y, AND2_38_Y, AND2_57_Y, 
        AO1_32_Y, AND2_3_Y, AO1_0_Y, AND2_53_Y, AND2_0_Y, AND2_60_Y, 
        AND2_34_Y, AND2_61_Y, AND2_12_Y, AND2_32_Y, AND2_26_Y, 
        AND2_36_Y, AND2_59_Y, AO1_30_Y, AND2_44_Y, AND2_58_Y, AO1_14_Y, 
        AO1_23_Y, AO1_6_Y, AO1_11_Y, AO1_2_Y, AO1_21_Y, AO1_18_Y, 
        AO1_7_Y, AO1_16_Y, AO1_35_Y, AO1_33_Y, XOR2_35_Y, XOR2_32_Y, 
        XOR2_47_Y, XOR2_69_Y, XOR2_18_Y, XOR2_63_Y, XOR2_58_Y, 
        XOR2_70_Y, XOR2_8_Y, XOR2_26_Y, XOR2_73_Y, XOR2_72_Y, 
        NAND2_1_Y, XOR2_28_Y, XOR2_24_Y, XOR2_15_Y, XOR2_49_Y, 
        XOR2_44_Y, XOR2_25_Y, XOR2_36_Y, XOR2_42_Y, XOR2_43_Y, 
        XOR2_13_Y, XOR2_37_Y, XOR2_1_Y, AND2_42_Y, AND2_9_Y, AND2_6_Y, 
        AND2_46_Y, AND2_10_Y, AND2_49_Y, AND2_14_Y, AND2_55_Y, 
        AND2_47_Y, AND2_2_Y, AND2_5_Y, XOR2_34_Y, XOR2_27_Y, XOR2_14_Y, 
        XOR2_61_Y, XOR2_57_Y, XOR2_54_Y, XOR2_0_Y, XOR2_45_Y, 
        XOR2_17_Y, XOR2_39_Y, XOR2_56_Y, XOR2_21_Y, AND2_11_Y, 
        AO1_20_Y, AND2_52_Y, AO1_3_Y, AND2_51_Y, AO1_4_Y, AND2_56_Y, 
        AO1_17_Y, AND2_41_Y, AO1_34_Y, AND2_8_Y, AND2_13_Y, AO1_22_Y, 
        AND2_27_Y, AO1_27_Y, AND2_23_Y, AND2_40_Y, AO1_13_Y, AND2_37_Y, 
        AND2_20_Y, AND2_19_Y, AND2_21_Y, AND2_7_Y, AND2_35_Y, 
        AND2_39_Y, AND2_48_Y, AND2_25_Y, AO1_1_Y, AO1_25_Y, AO1_24_Y, 
        AO1_19_Y, AO1_9_Y, AO1_10_Y, AO1_5_Y, AO1_26_Y, AO1_12_Y, 
        AO1_28_Y, XOR2_65_Y, XOR2_52_Y, XOR2_55_Y, XOR2_19_Y, 
        XOR2_33_Y, XOR2_7_Y, XOR2_64_Y, XOR2_71_Y, XOR2_31_Y, 
        XOR2_22_Y, XOR2_66_Y, \RAM4K9_QXI[0]_DOUTA0 , 
        \RAM4K9_QXI[1]_DOUTA0 , \RAM4K9_QXI[2]_DOUTA0 , 
        \RAM4K9_QXI[3]_DOUTA0 , \RAM4K9_QXI[4]_DOUTA0 , 
        \RAM4K9_QXI[5]_DOUTA0 , \RAM4K9_QXI[6]_DOUTA0 , 
        \RAM4K9_QXI[7]_DOUTA0 , \RAM4K9_QXI[0]_DOUTA1 , 
        \RAM4K9_QXI[1]_DOUTA1 , \RAM4K9_QXI[2]_DOUTA1 , 
        \RAM4K9_QXI[3]_DOUTA1 , \RAM4K9_QXI[4]_DOUTA1 , 
        \RAM4K9_QXI[5]_DOUTA1 , \RAM4K9_QXI[6]_DOUTA1 , 
        \RAM4K9_QXI[7]_DOUTA1 , AND3_0_Y, XNOR2_20_Y, XNOR2_10_Y, 
        XNOR2_6_Y, XNOR2_11_Y, XNOR2_12_Y, XNOR2_22_Y, XNOR2_9_Y, 
        XNOR2_16_Y, XNOR2_18_Y, XNOR2_14_Y, XNOR2_8_Y, XNOR2_21_Y, 
        AND3_7_Y, AND3_8_Y, AND3_9_Y, AND3_6_Y, AND2A_0_Y, AND3_1_Y, 
        XOR2_38_Y, XNOR2_1_Y, XNOR2_15_Y, XNOR2_19_Y, XNOR2_17_Y, 
        XNOR2_0_Y, XNOR2_4_Y, XNOR2_13_Y, XNOR2_7_Y, XNOR2_2_Y, 
        XNOR2_3_Y, XNOR2_5_Y, AND3_5_Y, AND3_2_Y, AND3_4_Y, AND3_3_Y, 
        NAND2_0_Y, VCC, GND;
    wire GND_power_net1;
    wire VCC_power_net1;
    assign GND = GND_power_net1;
    assign VCC = VCC_power_net1;
    
    AND2 AND2_2 (.A(\WBINSYNCSHIFT[11] ), .B(GND), .Y(AND2_2_Y));
    AND3 AND3_6 (.A(XNOR2_12_Y), .B(XNOR2_22_Y), .C(XNOR2_9_Y), .Y(
        AND3_6_Y));
    AND2 AND2_20 (.A(AND2_13_Y), .B(AND2_51_Y), .Y(AND2_20_Y));
    XNOR2 XNOR2_13 (.A(\MEM_RADDR[7] ), .B(\WBINNXTSHIFT[6] ), .Y(
        XNOR2_13_Y));
    AO1 AO1_11 (.A(XOR2_10_Y), .B(AO1_6_Y), .C(AND2_4_Y), .Y(AO1_11_Y));
    AND2 AND2_11 (.A(XOR2_34_Y), .B(XOR2_27_Y), .Y(AND2_11_Y));
    XOR2 \XOR2_WBINNXTSHIFT[2]  (.A(XOR2_52_Y), .B(AO1_1_Y), .Y(
        \WBINNXTSHIFT[2] ));
    AND2 AND2_22 (.A(\MEM_RADDR[8] ), .B(GND), .Y(AND2_22_Y));
    DFN1C0 \DFN1C0_RGRY[9]  (.D(XOR2_29_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[9] ));
    DFN1C0 DFN1C0_FULL (.D(FULLINT), .CLK(CLK), .CLR(READ_RESET_P), .Q(
        FULL));
    XNOR2 XNOR2_9 (.A(\RBINNXTSHIFT[6] ), .B(\WBINSYNCSHIFT[6] ), .Y(
        XNOR2_9_Y));
    XOR2 XOR2_19 (.A(\WBINSYNCSHIFT[5] ), .B(GND), .Y(XOR2_19_Y));
    AND2 AND2_44 (.A(AND2_60_Y), .B(XOR2_68_Y), .Y(AND2_44_Y));
    RAM4K9 \RAM4K9_QXI[6]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[14]), 
        .DINA0(DATA[6]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[6]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[6]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[6] ));
    AO1 AO1_31 (.A(XOR2_60_Y), .B(AND2_22_Y), .C(AND2_31_Y), .Y(
        AO1_31_Y));
    XOR2 XOR2_1 (.A(\WBINNXTSHIFT[11] ), .B(GND), .Y(XOR2_1_Y));
    XOR2 XOR2_23 (.A(\MEM_RADDR[5] ), .B(GND), .Y(XOR2_23_Y));
    DFN1E1C0 \DFN1E1C0_Q[1]  (.D(\QXI[1] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[1]));
    DFN1E1C0 \DFN1E1C0_Q[4]  (.D(\QXI[4] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[4]));
    DFN1E1C0 \DFN1E1C0_Q[7]  (.D(\QXI[7] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[7]));
    XOR2 XOR2_47 (.A(\MEM_RADDR[3] ), .B(GND), .Y(XOR2_47_Y));
    XOR2 XOR2_38 (.A(\MEM_RADDR[12] ), .B(\WBINNXTSHIFT[11] ), .Y(
        XOR2_38_Y));
    XOR2 \XOR2_RBINNXTSHIFT[0]  (.A(\MEM_RADDR[0] ), .B(MEMORYRE), .Y(
        \RBINNXTSHIFT[0] ));
    AO1 AO1_7 (.A(XOR2_12_Y), .B(AO1_18_Y), .C(AND2_22_Y), .Y(AO1_7_Y));
    DFN1C0 \DFN1C0_WGRY[6]  (.D(XOR2_36_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[6] ));
    AND2 AND2_18 (.A(XOR2_10_Y), .B(XOR2_23_Y), .Y(AND2_18_Y));
    AND2 AND2_15 (.A(\MEM_RADDR[5] ), .B(GND), .Y(AND2_15_Y));
    AO1 AO1_25 (.A(XOR2_14_Y), .B(AO1_1_Y), .C(AND2_9_Y), .Y(AO1_25_Y));
    XOR2 XOR2_45 (.A(\WBINSYNCSHIFT[8] ), .B(GND), .Y(XOR2_45_Y));
    XOR2 \XOR2_RBINNXTSHIFT[9]  (.A(XOR2_8_Y), .B(AO1_7_Y), .Y(
        \RBINNXTSHIFT[9] ));
    AND2 AND2_1 (.A(\MEM_RADDR[6] ), .B(GND), .Y(AND2_1_Y));
    XNOR2 XNOR2_21 (.A(\RBINNXTSHIFT[11] ), .B(\WBINSYNCSHIFT[11] ), 
        .Y(XNOR2_21_Y));
    AND2 AND2_49 (.A(\WBINSYNCSHIFT[7] ), .B(GND), .Y(AND2_49_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[1]  (.D(\RBINNXTSHIFT[1] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[1] ));
    AO1 AO1_8 (.A(XOR2_23_Y), .B(AND2_4_Y), .C(AND2_15_Y), .Y(AO1_8_Y));
    AND2 AND2_10 (.A(\WBINSYNCSHIFT[6] ), .B(GND), .Y(AND2_10_Y));
    AND2 AND2_7 (.A(AND2_13_Y), .B(XOR2_57_Y), .Y(AND2_7_Y));
    XOR2 XOR2_20 (.A(\RBINNXTSHIFT[1] ), .B(\RBINNXTSHIFT[2] ), .Y(
        XOR2_20_Y));
    XOR2 XOR2_63 (.A(\MEM_RADDR[6] ), .B(GND), .Y(XOR2_63_Y));
    RAM4K9 \RAM4K9_QXI[2]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[10]), 
        .DINA0(DATA[2]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[2]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[2]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[2] ));
    AND2 AND2_12 (.A(AND2_17_Y), .B(XOR2_9_Y), .Y(AND2_12_Y));
    DFN1C0 \DFN1C0_WGRY[5]  (.D(XOR2_25_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[5] ));
    XOR2 XOR2_52 (.A(\WBINSYNCSHIFT[3] ), .B(GND), .Y(XOR2_52_Y));
    AND2 AND2_61 (.A(AND2_0_Y), .B(AND2_45_Y), .Y(AND2_61_Y));
    AO1 AO1_15 (.A(XOR2_6_Y), .B(AND2_24_Y), .C(AND2_30_Y), .Y(
        AO1_15_Y));
    XOR2 \XOR2_WBINNXTSHIFT[0]  (.A(\WBINSYNCSHIFT[1] ), .B(MEMORYWE), 
        .Y(\WBINNXTSHIFT[0] ));
    DFN1C0 \DFN1C0_WGRY[7]  (.D(XOR2_42_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[7] ));
    AND2 AND2_EMPTYINT (.A(AND3_0_Y), .B(XNOR2_20_Y), .Y(EMPTYINT));
    XOR2 XOR2_24 (.A(\WBINNXTSHIFT[1] ), .B(\WBINNXTSHIFT[2] ), .Y(
        XOR2_24_Y));
    AND2 AND2_57 (.A(AND2_17_Y), .B(AND2_50_Y), .Y(AND2_57_Y));
    XOR2 XOR2_21 (.A(\WBINSYNCSHIFT[12] ), .B(GND), .Y(XOR2_21_Y));
    AO1 AO1_35 (.A(XOR2_46_Y), .B(AO1_16_Y), .C(AND2_24_Y), .Y(
        AO1_35_Y));
    XOR2 \XOR2_WBINNXTSHIFT[9]  (.A(XOR2_31_Y), .B(AO1_26_Y), .Y(
        \WBINNXTSHIFT[9] ));
    AND2 AND2_46 (.A(\WBINSYNCSHIFT[5] ), .B(GND), .Y(AND2_46_Y));
    XOR2 \XOR2_RBINNXTSHIFT[8]  (.A(XOR2_70_Y), .B(AO1_18_Y), .Y(
        \RBINNXTSHIFT[8] ));
    XOR2 XOR2_16 (.A(\RBINNXTSHIFT[7] ), .B(\RBINNXTSHIFT[8] ), .Y(
        XOR2_16_Y));
    XOR2 XOR2_60 (.A(\MEM_RADDR[9] ), .B(GND), .Y(XOR2_60_Y));
    AND2 AND2_43 (.A(\MEM_RADDR[3] ), .B(GND), .Y(AND2_43_Y));
    AO1 AO1_24 (.A(AND2_52_Y), .B(AO1_1_Y), .C(AO1_20_Y), .Y(AO1_24_Y));
    AND3 AND3_3 (.A(XNOR2_17_Y), .B(XNOR2_0_Y), .C(XNOR2_4_Y), .Y(
        AND3_3_Y));
    INV MEMWEBUBBLE (.A(MEMORYWE), .Y(MEMWENEG));
    AND2 AND2_6 (.A(\WBINSYNCSHIFT[4] ), .B(GND), .Y(AND2_6_Y));
    XOR2 XOR2_64 (.A(\WBINSYNCSHIFT[8] ), .B(GND), .Y(XOR2_64_Y));
    RAM4K9 \RAM4K9_QXI[1]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[9]), 
        .DINA0(DATA[1]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[1]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[1]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[1] ));
    AND3 AND3_0 (.A(AND3_8_Y), .B(XNOR2_8_Y), .C(XNOR2_21_Y), .Y(
        AND3_0_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[2]  (.D(\RBINNXTSHIFT[2] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[2] ));
    AND2 AND2_60 (.A(AND2_0_Y), .B(AND2_53_Y), .Y(AND2_60_Y));
    XOR2 XOR2_61 (.A(\WBINSYNCSHIFT[4] ), .B(GND), .Y(XOR2_61_Y));
    XOR2 XOR2_57 (.A(\WBINSYNCSHIFT[5] ), .B(GND), .Y(XOR2_57_Y));
    DFN1C0 \DFN1C0_RGRY[2]  (.D(XOR2_40_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[2] ));
    XOR2 XOR2_33 (.A(\WBINSYNCSHIFT[6] ), .B(GND), .Y(XOR2_33_Y));
    XNOR2 XNOR2_2 (.A(\MEM_RADDR[9] ), .B(\WBINNXTSHIFT[8] ), .Y(
        XNOR2_2_Y));
    XNOR2 XNOR2_19 (.A(\MEM_RADDR[3] ), .B(\WBINNXTSHIFT[2] ), .Y(
        XNOR2_19_Y));
    XOR2 XOR2_49 (.A(\WBINNXTSHIFT[3] ), .B(\WBINNXTSHIFT[4] ), .Y(
        XOR2_49_Y));
    XOR2 \XOR2_WBINNXTSHIFT[8]  (.A(XOR2_71_Y), .B(AO1_5_Y), .Y(
        \WBINNXTSHIFT[8] ));
    AO1 AO1_14 (.A(XOR2_5_Y), .B(AND2_58_Y), .C(AND2_33_Y), .Y(
        AO1_14_Y));
    XOR2 XOR2_4 (.A(\RBINNXTSHIFT[11] ), .B(\RBINNXTSHIFT[12] ), .Y(
        XOR2_4_Y));
    AND3 AND3_1 (.A(AND3_2_Y), .B(XNOR2_3_Y), .C(XNOR2_5_Y), .Y(
        AND3_1_Y));
    XOR2 XOR2_55 (.A(\WBINSYNCSHIFT[4] ), .B(GND), .Y(XOR2_55_Y));
    AND2 AND2_24 (.A(\MEM_RADDR[10] ), .B(GND), .Y(AND2_24_Y));
    XOR2 XOR2_72 (.A(\MEM_RADDR[12] ), .B(GND), .Y(XOR2_72_Y));
    XNOR2 XNOR2_0 (.A(\MEM_RADDR[5] ), .B(\WBINNXTSHIFT[4] ), .Y(
        XNOR2_0_Y));
    AND2 AND2_31 (.A(\MEM_RADDR[9] ), .B(GND), .Y(AND2_31_Y));
    AO1 AO1_34 (.A(XOR2_21_Y), .B(AND2_2_Y), .C(AND2_5_Y), .Y(AO1_34_Y)
        );
    XOR2 \XOR2_RBINNXTSHIFT[12]  (.A(XOR2_72_Y), .B(AO1_33_Y), .Y(
        \RBINNXTSHIFT[12] ));
    XOR2 XOR2_18 (.A(\MEM_RADDR[5] ), .B(GND), .Y(XOR2_18_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[2]  (.D(\WBINNXTSHIFT[1] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[2] ));
    DFN1C0 \DFN1C0_RGRY[11]  (.D(XOR2_4_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[11] ));
    XOR2 \XOR2_RBINNXTSHIFT[4]  (.A(XOR2_69_Y), .B(AO1_6_Y), .Y(
        \RBINNXTSHIFT[4] ));
    DFN1C0 \DFN1C0_RGRY[1]  (.D(XOR2_20_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[1] ));
    DFN1C0 \DFN1C0_WGRY[3]  (.D(XOR2_49_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[3] ));
    XOR2 XOR2_8 (.A(\MEM_RADDR[9] ), .B(GND), .Y(XOR2_8_Y));
    DFN1E1C0 \DFN1E1C0_Q[6]  (.D(\QXI[6] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[6]));
    XOR2 \XOR2_RBINNXTSHIFT[6]  (.A(XOR2_63_Y), .B(AO1_2_Y), .Y(
        \RBINNXTSHIFT[6] ));
    XOR2 XOR2_30 (.A(\RBINNXTSHIFT[12] ), .B(GND), .Y(XOR2_30_Y));
    AND2 AND2_38 (.A(XOR2_46_Y), .B(XOR2_6_Y), .Y(AND2_38_Y));
    AND2 AND2_35 (.A(AND2_20_Y), .B(XOR2_0_Y), .Y(AND2_35_Y));
    INV MEMREBUBBLE (.A(MEMORYRE), .Y(MEMRENEG));
    DFN1C0 \DFN1C0_WGRY[11]  (.D(XOR2_1_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[11] ));
    AND2 AND2_29 (.A(XOR2_48_Y), .B(XOR2_3_Y), .Y(AND2_29_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[4]  (.D(\RBINNXTSHIFT[4] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[4] ));
    XOR2 XOR2_34 (.A(\WBINSYNCSHIFT[1] ), .B(MEMORYWE), .Y(XOR2_34_Y));
    XOR2 XOR2_31 (.A(\WBINSYNCSHIFT[10] ), .B(GND), .Y(XOR2_31_Y));
    AND2 AND2_3 (.A(AND2_18_Y), .B(AND2_29_Y), .Y(AND2_3_Y));
    AND2 AND2_30 (.A(\MEM_RADDR[11] ), .B(GND), .Y(AND2_30_Y));
    XOR2 \XOR2_WBINNXTSHIFT[4]  (.A(XOR2_19_Y), .B(AO1_24_Y), .Y(
        \WBINNXTSHIFT[4] ));
    XNOR2 XNOR2_6 (.A(\RBINNXTSHIFT[2] ), .B(\WBINSYNCSHIFT[2] ), .Y(
        XNOR2_6_Y));
    AND2 AND2_14 (.A(\WBINSYNCSHIFT[8] ), .B(GND), .Y(AND2_14_Y));
    INV RESETBUBBLE (.A(RESET), .Y(READ_RESET_P));
    AND2 AND2_32 (.A(AND2_57_Y), .B(XOR2_10_Y), .Y(AND2_32_Y));
    XOR2 \XOR2_WBINNXTSHIFT[6]  (.A(XOR2_7_Y), .B(AO1_9_Y), .Y(
        \WBINNXTSHIFT[6] ));
    DFN1C0 \DFN1C0_MEM_RADDR[5]  (.D(\RBINNXTSHIFT[5] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[5] ));
    AND3 AND3_8 (.A(AND3_9_Y), .B(AND3_7_Y), .C(AND3_6_Y), .Y(AND3_8_Y)
        );
    XOR2 XOR2_46 (.A(\MEM_RADDR[10] ), .B(GND), .Y(XOR2_46_Y));
    XNOR2 XNOR2_11 (.A(\RBINNXTSHIFT[3] ), .B(\WBINSYNCSHIFT[3] ), .Y(
        XNOR2_11_Y));
    AO1 AO1_2 (.A(AND2_18_Y), .B(AO1_6_Y), .C(AO1_8_Y), .Y(AO1_2_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[8]  (.D(\RBINNXTSHIFT[8] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[8] ));
    DFN1C0 \DFN1C0_WGRY[0]  (.D(XOR2_28_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[0] ));
    AND2 AND2_26 (.A(AND2_34_Y), .B(XOR2_48_Y), .Y(AND2_26_Y));
    RAM4K9 \RAM4K9_QXI[7]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[15]), 
        .DINA0(DATA[7]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[7]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[7]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[7] ));
    XOR2 XOR2_9 (.A(\MEM_RADDR[2] ), .B(GND), .Y(XOR2_9_Y));
    AND3 AND3_5 (.A(XNOR2_1_Y), .B(XNOR2_15_Y), .C(XNOR2_19_Y), .Y(
        AND3_5_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[1]  (.D(\WBINNXTSHIFT[0] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[1] ));
    XOR2 XOR2_59 (.A(\RBINNXTSHIFT[4] ), .B(\RBINNXTSHIFT[5] ), .Y(
        XOR2_59_Y));
    AND2 AND2_23 (.A(AND2_41_Y), .B(AND2_8_Y), .Y(AND2_23_Y));
    XNOR2 XNOR2_4 (.A(\MEM_RADDR[6] ), .B(\WBINNXTSHIFT[5] ), .Y(
        XNOR2_4_Y));
    DFN1C0 \DFN1C0_RGRY[8]  (.D(XOR2_50_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[8] ));
    XOR2 XOR2_5 (.A(\MEM_RADDR[1] ), .B(GND), .Y(XOR2_5_Y));
    XNOR2 XNOR2_20 (.A(\RBINNXTSHIFT[12] ), .B(\WBINSYNCSHIFT[12] ), 
        .Y(XNOR2_20_Y));
    AO1 AO1_28 (.A(XOR2_56_Y), .B(AO1_12_Y), .C(AND2_2_Y), .Y(AO1_28_Y)
        );
    AND2 AND2_19 (.A(AND2_40_Y), .B(AND2_41_Y), .Y(AND2_19_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[6]  (.D(\RBINNXTSHIFT[6] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[6] ));
    DFN1E1C0 \DFN1E1C0_Q[0]  (.D(\QXI[0] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[0]));
    XOR2 XOR2_22 (.A(\WBINSYNCSHIFT[11] ), .B(GND), .Y(XOR2_22_Y));
    AO1 AO1_1 (.A(XOR2_27_Y), .B(AND2_25_Y), .C(AND2_42_Y), .Y(AO1_1_Y)
        );
    XOR2 XOR2_13 (.A(\WBINNXTSHIFT[9] ), .B(\WBINNXTSHIFT[10] ), .Y(
        XOR2_13_Y));
    XNOR2 XNOR2_18 (.A(\RBINNXTSHIFT[8] ), .B(\WBINSYNCSHIFT[8] ), .Y(
        XNOR2_18_Y));
    AND2 AND2_51 (.A(XOR2_57_Y), .B(XOR2_54_Y), .Y(AND2_51_Y));
    AO1 AO1_3 (.A(XOR2_54_Y), .B(AND2_46_Y), .C(AND2_10_Y), .Y(AO1_3_Y)
        );
    AND2 AND2_47 (.A(\WBINSYNCSHIFT[10] ), .B(GND), .Y(AND2_47_Y));
    AO1 AO1_18 (.A(AND2_3_Y), .B(AO1_6_Y), .C(AO1_32_Y), .Y(AO1_18_Y));
    XOR2 XOR2_48 (.A(\MEM_RADDR[6] ), .B(GND), .Y(XOR2_48_Y));
    XOR2 \XOR2_RBINNXTSHIFT[3]  (.A(XOR2_47_Y), .B(AO1_23_Y), .Y(
        \RBINNXTSHIFT[3] ));
    DFN1C0 \DFN1C0_MEM_RADDR[7]  (.D(\RBINNXTSHIFT[7] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[7] ));
    AND2 AND2_16 (.A(\MEM_RADDR[2] ), .B(GND), .Y(AND2_16_Y));
    DFN1C0 \DFN1C0_WGRY[9]  (.D(XOR2_13_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[9] ));
    XOR2 XOR2_62 (.A(\RBINNXTSHIFT[10] ), .B(\RBINNXTSHIFT[11] ), .Y(
        XOR2_62_Y));
    AND2 AND2_13 (.A(AND2_11_Y), .B(AND2_52_Y), .Y(AND2_13_Y));
    XOR2 XOR2_10 (.A(\MEM_RADDR[4] ), .B(GND), .Y(XOR2_10_Y));
    XNOR2 XNOR2_1 (.A(\MEM_RADDR[1] ), .B(\WBINNXTSHIFT[0] ), .Y(
        XNOR2_1_Y));
    AND2 AND2_58 (.A(\MEM_RADDR[0] ), .B(MEMORYRE), .Y(AND2_58_Y));
    AND2 AND2_55 (.A(\WBINSYNCSHIFT[9] ), .B(GND), .Y(AND2_55_Y));
    RAM4K9 \RAM4K9_QXI[0]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[8]), 
        .DINA0(DATA[0]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[0]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[0]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[0] ));
    DFN1C0 \DFN1C0_RGRY[4]  (.D(XOR2_59_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[4] ));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[6]  (.D(\WBINNXTSHIFT[5] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[6] ));
    XOR2 XOR2_27 (.A(\WBINSYNCSHIFT[2] ), .B(GND), .Y(XOR2_27_Y));
    AND2 AND2_MEMORYRE (.A(NAND2_1_Y), .B(RE), .Y(MEMORYRE));
    XOR2 \XOR2_WBINNXTSHIFT[3]  (.A(XOR2_55_Y), .B(AO1_25_Y), .Y(
        \WBINNXTSHIFT[3] ));
    XOR2 XOR2_7 (.A(\WBINSYNCSHIFT[7] ), .B(GND), .Y(XOR2_7_Y));
    AND2 AND2_5 (.A(\WBINSYNCSHIFT[12] ), .B(GND), .Y(AND2_5_Y));
    XOR2 XOR2_56 (.A(\WBINSYNCSHIFT[11] ), .B(GND), .Y(XOR2_56_Y));
    RAM4K9 \RAM4K9_QXI[4]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[12]), 
        .DINA0(DATA[4]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[4]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[4]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[4] ));
    XOR2 XOR2_14 (.A(\WBINSYNCSHIFT[3] ), .B(GND), .Y(XOR2_14_Y));
    AND2 AND2_50 (.A(XOR2_9_Y), .B(XOR2_2_Y), .Y(AND2_50_Y));
    XNOR2 XNOR2_3 (.A(\MEM_RADDR[10] ), .B(\WBINNXTSHIFT[9] ), .Y(
        XNOR2_3_Y));
    XOR2 XOR2_11 (.A(\RBINNXTSHIFT[0] ), .B(\RBINNXTSHIFT[1] ), .Y(
        XOR2_11_Y));
    XNOR2 XNOR2_22 (.A(\RBINNXTSHIFT[5] ), .B(\WBINSYNCSHIFT[5] ), .Y(
        XNOR2_22_Y));
    AND2 AND2_52 (.A(XOR2_14_Y), .B(XOR2_61_Y), .Y(AND2_52_Y));
    XOR2 XOR2_25 (.A(\WBINNXTSHIFT[5] ), .B(\WBINNXTSHIFT[6] ), .Y(
        XOR2_25_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[4]  (.D(\WBINNXTSHIFT[3] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[4] ));
    XNOR2 XNOR2_15 (.A(\MEM_RADDR[2] ), .B(\WBINNXTSHIFT[1] ), .Y(
        XNOR2_15_Y));
    AO1 AO1_22 (.A(AND2_56_Y), .B(AO1_3_Y), .C(AO1_4_Y), .Y(AO1_22_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[12]  (.D(\WBINNXTSHIFT[11] ), .CLK(
        CLK), .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[12] ));
    AND2 AND2_34 (.A(AND2_57_Y), .B(AND2_18_Y), .Y(AND2_34_Y));
    AO1 AO1_6 (.A(AND2_50_Y), .B(AO1_14_Y), .C(AO1_29_Y), .Y(AO1_6_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[3]  (.D(\RBINNXTSHIFT[3] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[3] ));
    XOR2 XOR2_67 (.A(\RBINNXTSHIFT[5] ), .B(\RBINNXTSHIFT[6] ), .Y(
        XOR2_67_Y));
    AND3 AND3_2 (.A(AND3_4_Y), .B(AND3_5_Y), .C(AND3_3_Y), .Y(AND3_2_Y)
        );
    AO1 AO1_12 (.A(AND2_41_Y), .B(AO1_5_Y), .C(AO1_17_Y), .Y(AO1_12_Y));
    XOR2 XOR2_32 (.A(\MEM_RADDR[2] ), .B(GND), .Y(XOR2_32_Y));
    AND2 AND2_9 (.A(\WBINSYNCSHIFT[3] ), .B(GND), .Y(AND2_9_Y));
    DFN1E1C0 \DFN1E1C0_Q[5]  (.D(\QXI[5] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[5]));
    XOR2 XOR2_65 (.A(\WBINSYNCSHIFT[2] ), .B(GND), .Y(XOR2_65_Y));
    XOR2 XOR2_58 (.A(\MEM_RADDR[7] ), .B(GND), .Y(XOR2_58_Y));
    AO1 AO1_32 (.A(AND2_29_Y), .B(AO1_8_Y), .C(AO1_36_Y), .Y(AO1_32_Y));
    XOR2 XOR2_43 (.A(\WBINNXTSHIFT[8] ), .B(\WBINNXTSHIFT[9] ), .Y(
        XOR2_43_Y));
    AO1 AO1_9 (.A(AND2_51_Y), .B(AO1_24_Y), .C(AO1_3_Y), .Y(AO1_9_Y));
    DFN1C0 DFN1C0_DVLDX (.D(DVLDI), .CLK(CLK), .CLR(READ_RESET_P), .Q(
        DVLDX));
    AND2 AND2_39 (.A(AND2_40_Y), .B(XOR2_17_Y), .Y(AND2_39_Y));
    NAND2 NAND2_0 (.A(FULL), .B(VCC), .Y(NAND2_0_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[7]  (.D(\WBINNXTSHIFT[6] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[7] ));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[11]  (.D(\WBINNXTSHIFT[10] ), .CLK(
        CLK), .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[11] ));
    DFN1C0 \DFN1C0_RGRY[6]  (.D(XOR2_51_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[6] ));
    AND2 AND2_27 (.A(AND2_51_Y), .B(AND2_56_Y), .Y(AND2_27_Y));
    DFN1C0 DFN1C0_DVLDI (.D(AND2A_0_Y), .CLK(CLK), .CLR(READ_RESET_P), 
        .Q(DVLDI));
    XNOR2 XNOR2_10 (.A(\RBINNXTSHIFT[1] ), .B(\WBINSYNCSHIFT[1] ), .Y(
        XNOR2_10_Y));
    AND2 AND2_MEMORYWE (.A(NAND2_0_Y), .B(WE), .Y(MEMORYWE));
    AO1 AO1_20 (.A(XOR2_61_Y), .B(AND2_9_Y), .C(AND2_6_Y), .Y(AO1_20_Y)
        );
    DFN1C0 \DFN1C0_WGRY[2]  (.D(XOR2_15_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[2] ));
    AO1 AO1_0 (.A(AND2_38_Y), .B(AO1_31_Y), .C(AO1_15_Y), .Y(AO1_0_Y));
    XOR2 XOR2_29 (.A(\RBINNXTSHIFT[9] ), .B(\RBINNXTSHIFT[10] ), .Y(
        XOR2_29_Y));
    XOR2 XOR2_40 (.A(\RBINNXTSHIFT[2] ), .B(\RBINNXTSHIFT[3] ), .Y(
        XOR2_40_Y));
    XOR2 XOR2_2 (.A(\MEM_RADDR[3] ), .B(GND), .Y(XOR2_2_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[9]  (.D(\WBINNXTSHIFT[8] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[9] ));
    DFN1C0 \DFN1C0_RGRY[5]  (.D(XOR2_67_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[5] ));
    AND2 AND2_36 (.A(AND2_0_Y), .B(XOR2_12_Y), .Y(AND2_36_Y));
    XOR2 XOR2_37 (.A(\WBINNXTSHIFT[10] ), .B(\WBINNXTSHIFT[11] ), .Y(
        XOR2_37_Y));
    AND2A AND2A_0 (.A(EMPTY), .B(RE), .Y(AND2A_0_Y));
    AO1 AO1_26 (.A(XOR2_17_Y), .B(AO1_5_Y), .C(AND2_55_Y), .Y(AO1_26_Y)
        );
    DFN1C0 \DFN1C0_WGRY[10]  (.D(XOR2_37_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[10] ));
    DFN1C0 \DFN1C0_RGRY[7]  (.D(XOR2_16_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[7] ));
    AND3 AND3_9 (.A(XNOR2_16_Y), .B(XNOR2_18_Y), .C(XNOR2_14_Y), .Y(
        AND3_9_Y));
    XOR2 \XOR2_RBINNXTSHIFT[5]  (.A(XOR2_18_Y), .B(AO1_11_Y), .Y(
        \RBINNXTSHIFT[5] ));
    AO1 AO1_23 (.A(XOR2_9_Y), .B(AO1_14_Y), .C(AND2_16_Y), .Y(AO1_23_Y)
        );
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[3]  (.D(\WBINNXTSHIFT[2] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[3] ));
    AND2 AND2_33 (.A(\MEM_RADDR[1] ), .B(GND), .Y(AND2_33_Y));
    XOR2 XOR2_44 (.A(\WBINNXTSHIFT[4] ), .B(\WBINNXTSHIFT[5] ), .Y(
        XOR2_44_Y));
    AO1 AO1_10 (.A(XOR2_0_Y), .B(AO1_9_Y), .C(AND2_49_Y), .Y(AO1_10_Y));
    XOR2 XOR2_41 (.A(\RBINNXTSHIFT[3] ), .B(\RBINNXTSHIFT[4] ), .Y(
        XOR2_41_Y));
    XOR2 XOR2_35 (.A(\MEM_RADDR[1] ), .B(GND), .Y(XOR2_35_Y));
    XOR2 \XOR2_RBINNXTSHIFT[10]  (.A(XOR2_26_Y), .B(AO1_16_Y), .Y(
        \RBINNXTSHIFT[10] ));
    DFN1C0 \DFN1C0_WGRY[1]  (.D(XOR2_24_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[1] ));
    DFN1P0 DFN1P0_EMPTY (.D(EMPTYINT), .CLK(CLK), .PRE(READ_RESET_P), 
        .Q(EMPTY));
    DFN1E1C0 \DFN1E1C0_Q[3]  (.D(\QXI[3] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[3]));
    AO1 AO1_30 (.A(XOR2_68_Y), .B(AO1_33_Y), .C(AND2_54_Y), .Y(
        AO1_30_Y));
    XOR2 \XOR2_RBINNXTSHIFT[7]  (.A(XOR2_58_Y), .B(AO1_21_Y), .Y(
        \RBINNXTSHIFT[7] ));
    AND2 AND2_41 (.A(XOR2_17_Y), .B(XOR2_39_Y), .Y(AND2_41_Y));
    AND2 AND2_0 (.A(AND2_57_Y), .B(AND2_3_Y), .Y(AND2_0_Y));
    XOR2 XOR2_69 (.A(\MEM_RADDR[4] ), .B(GND), .Y(XOR2_69_Y));
    DFN1C0 \DFN1C0_RGRY[12]  (.D(XOR2_30_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[12] ));
    AO1 AO1_16 (.A(AND2_45_Y), .B(AO1_18_Y), .C(AO1_31_Y), .Y(AO1_16_Y)
        );
    AND2 AND2_17 (.A(XOR2_53_Y), .B(XOR2_5_Y), .Y(AND2_17_Y));
    AO1 AO1_29 (.A(XOR2_2_Y), .B(AND2_16_Y), .C(AND2_43_Y), .Y(
        AO1_29_Y));
    XOR2 XOR2_6 (.A(\MEM_RADDR[11] ), .B(GND), .Y(XOR2_6_Y));
    AND2 AND2_54 (.A(\MEM_RADDR[12] ), .B(GND), .Y(AND2_54_Y));
    AO1 AO1_13 (.A(AND2_23_Y), .B(AO1_5_Y), .C(AO1_27_Y), .Y(AO1_13_Y));
    XOR2 \XOR2_WBINNXTSHIFT[5]  (.A(XOR2_33_Y), .B(AO1_19_Y), .Y(
        \WBINNXTSHIFT[5] ));
    AO1 AO1_36 (.A(XOR2_3_Y), .B(AND2_1_Y), .C(AND2_28_Y), .Y(AO1_36_Y)
        );
    XOR2 XOR2_53 (.A(\MEM_RADDR[0] ), .B(MEMORYRE), .Y(XOR2_53_Y));
    AO1 AO1_33 (.A(AND2_53_Y), .B(AO1_18_Y), .C(AO1_0_Y), .Y(AO1_33_Y));
    XOR2 \XOR2_WBINNXTSHIFT[10]  (.A(XOR2_22_Y), .B(AO1_12_Y), .Y(
        \WBINNXTSHIFT[10] ));
    XNOR2 XNOR2_12 (.A(\RBINNXTSHIFT[4] ), .B(\WBINSYNCSHIFT[4] ), .Y(
        XNOR2_12_Y));
    XOR2 XOR2_12 (.A(\MEM_RADDR[8] ), .B(GND), .Y(XOR2_12_Y));
    XNOR2 XNOR2_7 (.A(\MEM_RADDR[8] ), .B(\WBINNXTSHIFT[7] ), .Y(
        XNOR2_7_Y));
    AND2 AND2_48 (.A(AND2_19_Y), .B(XOR2_56_Y), .Y(AND2_48_Y));
    AND2 AND2_45 (.A(XOR2_12_Y), .B(XOR2_60_Y), .Y(AND2_45_Y));
    AO1 AO1_19 (.A(XOR2_57_Y), .B(AO1_24_Y), .C(AND2_46_Y), .Y(
        AO1_19_Y));
    XOR2 \XOR2_WBINNXTSHIFT[7]  (.A(XOR2_64_Y), .B(AO1_10_Y), .Y(
        \WBINNXTSHIFT[7] ));
    RAM4K9 \RAM4K9_QXI[5]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[13]), 
        .DINA0(DATA[5]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[5]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[5]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[5] ));
    DFN1C0 \DFN1C0_MEM_RADDR[12]  (.D(\RBINNXTSHIFT[12] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[12] ));
    XOR2 XOR2_26 (.A(\MEM_RADDR[10] ), .B(GND), .Y(XOR2_26_Y));
    AND2 AND2_59 (.A(AND2_61_Y), .B(XOR2_46_Y), .Y(AND2_59_Y));
    DFN1C0 \DFN1C0_RGRY[10]  (.D(XOR2_62_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[10] ));
    AND2 AND2_4 (.A(\MEM_RADDR[4] ), .B(GND), .Y(AND2_4_Y));
    AND2 AND2_FULLINT (.A(AND3_1_Y), .B(XOR2_38_Y), .Y(FULLINT));
    AND2 AND2_40 (.A(AND2_13_Y), .B(AND2_27_Y), .Y(AND2_40_Y));
    XOR2 XOR2_50 (.A(\RBINNXTSHIFT[8] ), .B(\RBINNXTSHIFT[9] ), .Y(
        XOR2_50_Y));
    AND2 AND2_42 (.A(\WBINSYNCSHIFT[2] ), .B(GND), .Y(AND2_42_Y));
    DFN1E1C0 \DFN1E1C0_Q[2]  (.D(\QXI[2] ), .CLK(CLK), .CLR(
        READ_RESET_P), .E(DVLDI), .Q(Q[2]));
    DFN1C0 \DFN1C0_WGRY[8]  (.D(XOR2_43_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[8] ));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[8]  (.D(\WBINNXTSHIFT[7] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[8] ));
    XNOR2 XNOR2_5 (.A(\MEM_RADDR[11] ), .B(\WBINNXTSHIFT[10] ), .Y(
        XNOR2_5_Y));
    AO1 AO1_5 (.A(AND2_27_Y), .B(AO1_24_Y), .C(AO1_22_Y), .Y(AO1_5_Y));
    XNOR2 XNOR2_16 (.A(\RBINNXTSHIFT[7] ), .B(\WBINSYNCSHIFT[7] ), .Y(
        XNOR2_16_Y));
    DFN1C0 \DFN1C0_RGRY[3]  (.D(XOR2_41_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[3] ));
    XOR2 XOR2_39 (.A(\WBINSYNCSHIFT[10] ), .B(GND), .Y(XOR2_39_Y));
    AND2 AND2_8 (.A(XOR2_56_Y), .B(XOR2_21_Y), .Y(AND2_8_Y));
    XOR2 XOR2_3 (.A(\MEM_RADDR[7] ), .B(GND), .Y(XOR2_3_Y));
    XOR2 XOR2_54 (.A(\WBINSYNCSHIFT[6] ), .B(GND), .Y(XOR2_54_Y));
    XOR2 \XOR2_RBINNXTSHIFT[11]  (.A(XOR2_73_Y), .B(AO1_35_Y), .Y(
        \RBINNXTSHIFT[11] ));
    AO1 AO1_27 (.A(AND2_8_Y), .B(AO1_17_Y), .C(AO1_34_Y), .Y(AO1_27_Y));
    XOR2 XOR2_51 (.A(\RBINNXTSHIFT[6] ), .B(\RBINNXTSHIFT[7] ), .Y(
        XOR2_51_Y));
    XOR2 XOR2_66 (.A(\WBINSYNCSHIFT[12] ), .B(GND), .Y(XOR2_66_Y));
    AND2 AND2_56 (.A(XOR2_0_Y), .B(XOR2_45_Y), .Y(AND2_56_Y));
    XOR2 \XOR2_RBINNXTSHIFT[1]  (.A(XOR2_35_Y), .B(AND2_58_Y), .Y(
        \RBINNXTSHIFT[1] ));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[10]  (.D(\WBINNXTSHIFT[9] ), .CLK(CLK)
        , .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[10] ));
    XOR2 XOR2_17 (.A(\WBINSYNCSHIFT[9] ), .B(GND), .Y(XOR2_17_Y));
    XOR2 XOR2_73 (.A(\MEM_RADDR[11] ), .B(GND), .Y(XOR2_73_Y));
    AND2 AND2_53 (.A(AND2_45_Y), .B(AND2_38_Y), .Y(AND2_53_Y));
    AND3 AND3_7 (.A(XNOR2_10_Y), .B(XNOR2_6_Y), .C(XNOR2_11_Y), .Y(
        AND3_7_Y));
    XOR2 XOR2_28 (.A(\WBINNXTSHIFT[0] ), .B(\WBINNXTSHIFT[1] ), .Y(
        XOR2_28_Y));
    XOR2 XOR2_15 (.A(\WBINNXTSHIFT[2] ), .B(\WBINNXTSHIFT[3] ), .Y(
        XOR2_15_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[0]  (.D(\RBINNXTSHIFT[0] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[0] ));
    AO1 AO1_17 (.A(XOR2_39_Y), .B(AND2_55_Y), .C(AND2_47_Y), .Y(
        AO1_17_Y));
    XNOR2 XNOR2_17 (.A(\MEM_RADDR[4] ), .B(\WBINNXTSHIFT[3] ), .Y(
        XNOR2_17_Y));
    RAM4K9 \RAM4K9_QXI[3]  (.ADDRA11(GND), .ADDRA10(
        \WBINSYNCSHIFT[11] ), .ADDRA9(\WBINSYNCSHIFT[10] ), .ADDRA8(
        \WBINSYNCSHIFT[9] ), .ADDRA7(\WBINSYNCSHIFT[8] ), .ADDRA6(
        \WBINSYNCSHIFT[7] ), .ADDRA5(\WBINSYNCSHIFT[6] ), .ADDRA4(
        \WBINSYNCSHIFT[5] ), .ADDRA3(\WBINSYNCSHIFT[4] ), .ADDRA2(
        \WBINSYNCSHIFT[3] ), .ADDRA1(\WBINSYNCSHIFT[2] ), .ADDRA0(
        \WBINSYNCSHIFT[1] ), .ADDRB11(\MEM_RADDR[11] ), .ADDRB10(
        \MEM_RADDR[10] ), .ADDRB9(\MEM_RADDR[9] ), .ADDRB8(
        \MEM_RADDR[8] ), .ADDRB7(\MEM_RADDR[7] ), .ADDRB6(
        \MEM_RADDR[6] ), .ADDRB5(\MEM_RADDR[5] ), .ADDRB4(
        \MEM_RADDR[4] ), .ADDRB3(\MEM_RADDR[3] ), .ADDRB2(
        \MEM_RADDR[2] ), .ADDRB1(\MEM_RADDR[1] ), .ADDRB0(
        \MEM_RADDR[0] ), .DINA8(GND), .DINA7(GND), .DINA6(GND), .DINA5(
        GND), .DINA4(GND), .DINA3(GND), .DINA2(GND), .DINA1(DATA[11]), 
        .DINA0(DATA[3]), .DINB8(GND), .DINB7(GND), .DINB6(GND), .DINB5(
        GND), .DINB4(GND), .DINB3(GND), .DINB2(GND), .DINB1(GND), 
        .DINB0(GND), .WIDTHA0(VCC), .WIDTHA1(GND), .WIDTHB0(GND), 
        .WIDTHB1(GND), .PIPEA(GND), .PIPEB(GND), .WMODEA(GND), .WMODEB(
        GND), .BLKA(MEMWENEG), .BLKB(MEMRENEG), .WENA(GND), .WENB(VCC), 
        .CLKA(CLK), .CLKB(CLK), .RESET(READ_RESET_P), .DOUTA8(), 
        .DOUTA7(), .DOUTA6(), .DOUTA5(), .DOUTA4(), .DOUTA3(), .DOUTA2(
        ), .DOUTA1(\RAM4K9_QXI[3]_DOUTA1 ), .DOUTA0(
        \RAM4K9_QXI[3]_DOUTA0 ), .DOUTB8(), .DOUTB7(), .DOUTB6(), 
        .DOUTB5(), .DOUTB4(), .DOUTB3(), .DOUTB2(), .DOUTB1(), .DOUTB0(
        \QXI[3] ));
    DFN1C0 \DFN1C0_MEM_RADDR[10]  (.D(\RBINNXTSHIFT[10] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[10] ));
    XOR2 \XOR2_WBINNXTSHIFT[11]  (.A(XOR2_66_Y), .B(AO1_28_Y), .Y(
        \WBINNXTSHIFT[11] ));
    AND3 AND3_4 (.A(XNOR2_13_Y), .B(XNOR2_7_Y), .C(XNOR2_2_Y), .Y(
        AND3_4_Y));
    DFN1C0 \DFN1C0_RGRY[0]  (.D(XOR2_11_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\RGRY[0] ));
    XOR2 \XOR2_WBINNXTSHIFT[1]  (.A(XOR2_65_Y), .B(AND2_25_Y), .Y(
        \WBINNXTSHIFT[1] ));
    AND2 AND2_21 (.A(AND2_11_Y), .B(XOR2_14_Y), .Y(AND2_21_Y));
    DFN1C0 \DFN1C0_WGRY[4]  (.D(XOR2_44_Y), .CLK(CLK), .CLR(
        READ_RESET_P), .Q(\WGRY[4] ));
    XOR2 XOR2_0 (.A(\WBINSYNCSHIFT[7] ), .B(GND), .Y(XOR2_0_Y));
    XOR2 XOR2_70 (.A(\MEM_RADDR[8] ), .B(GND), .Y(XOR2_70_Y));
    NAND2 NAND2_1 (.A(EMPTY), .B(VCC), .Y(NAND2_1_Y));
    AO1 AO1_4 (.A(XOR2_45_Y), .B(AND2_49_Y), .C(AND2_14_Y), .Y(AO1_4_Y)
        );
    XOR2 XOR2_68 (.A(\MEM_RADDR[12] ), .B(GND), .Y(XOR2_68_Y));
    AND2 AND2_37 (.A(AND2_40_Y), .B(AND2_23_Y), .Y(AND2_37_Y));
    XNOR2 XNOR2_14 (.A(\RBINNXTSHIFT[9] ), .B(\WBINSYNCSHIFT[9] ), .Y(
        XNOR2_14_Y));
    XOR2 XOR2_42 (.A(\WBINNXTSHIFT[7] ), .B(\WBINNXTSHIFT[8] ), .Y(
        XOR2_42_Y));
    XOR2 \XOR2_RBINNXTSHIFT[2]  (.A(XOR2_32_Y), .B(AO1_14_Y), .Y(
        \RBINNXTSHIFT[2] ));
    AO1 AO1_21 (.A(XOR2_48_Y), .B(AO1_2_Y), .C(AND2_1_Y), .Y(AO1_21_Y));
    DFN1C0 \DFN1C0_MEM_RADDR[9]  (.D(\RBINNXTSHIFT[9] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[9] ));
    XOR2 XOR2_36 (.A(\WBINNXTSHIFT[6] ), .B(\WBINNXTSHIFT[7] ), .Y(
        XOR2_36_Y));
    XNOR2 XNOR2_8 (.A(\RBINNXTSHIFT[10] ), .B(\WBINSYNCSHIFT[10] ), .Y(
        XNOR2_8_Y));
    XOR2 XOR2_71 (.A(\WBINSYNCSHIFT[9] ), .B(GND), .Y(XOR2_71_Y));
    AND2 AND2_28 (.A(\MEM_RADDR[7] ), .B(GND), .Y(AND2_28_Y));
    AND2 AND2_25 (.A(\WBINSYNCSHIFT[1] ), .B(MEMORYWE), .Y(AND2_25_Y));
    DFN1C0 \DFN1C0_WBINSYNCSHIFT[5]  (.D(\WBINNXTSHIFT[4] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\WBINSYNCSHIFT[5] ));
    DFN1C0 \DFN1C0_MEM_RADDR[11]  (.D(\RBINNXTSHIFT[11] ), .CLK(CLK), 
        .CLR(READ_RESET_P), .Q(\MEM_RADDR[11] ));
    GND GND_power_inst1 (.Y(GND_power_net1));
    VCC VCC_power_inst1 (.Y(VCC_power_net1));
    
endmodule

// _Disclaimer: Please leave the following comments in the file, they are for internal purposes only._


// _GEN_File_Contents_

// Version:11.8.3.6
// ACTGENU_CALL:1
// BATCH:T
// FAM:PA3LC
// OUTFORMAT:Verilog
// LPMTYPE:LPM_SOFTFIFO
// LPM_HINT:MEMFF
// INSERT_PAD:NO
// INSERT_IOREG:NO
// GEN_BHV_VHDL_VAL:F
// GEN_BHV_VERILOG_VAL:F
// MGNTIMER:F
// MGNCMPL:T
// DESDIR:D:/NHI/fpga/top/MDM/Build_MDM/smartgen\FIFOCore_2Bto1B_2048
// GEN_BEHV_MODULE:F
// SMARTGEN_DIE:IS4X2M1
// SMARTGEN_PACKAGE:vq100
// AGENIII_IS_SUBPROJECT_LIBERO:T
// WWIDTH:16
// WDEPTH:2048
// RWIDTH:8
// RDEPTH:4096
// CLKS:1
// CLOCK_PN:CLK
// WCLK_EDGE:RISE
// ACLR_PN:RESET
// RESET_POLARITY:1
// INIT_RAM:F
// WE_POLARITY:1
// RE_POLARITY:1
// FF_PN:FULL
// AF_PN:AFULL
// WACK_PN:WACK
// OVRFLOW_PN:OVERFLOW
// WRCNT_PN:WRCNT
// WE_PN:WE
// EF_PN:EMPTY
// AE_PN:AEMPTY
// DVLD_PN:DVLD
// UDRFLOW_PN:UNDERFLOW
// RDCNT_PN:RDCNT
// RE_PN:RE
// CONTROLLERONLY:F
// FSTOP:YES
// ESTOP:YES
// WRITEACK:NO
// OVERFLOW:NO
// WRCOUNT:NO
// DATAVALID:NO
// UNDERFLOW:NO
// RDCOUNT:NO
// AF_PORT_PN:AFVAL
// AE_PORT_PN:AEVAL
// AFFLAG:NONE
// AEFLAG:NONE
// DATA_IN_PN:DATA
// DATA_OUT_PN:Q
// CASCADE:0

// _End_Comments_

